module wobbl_e_character_render(
	input[7:0] character,
	input[2:0] line_no,
	out[4:0] bit_row);
	

	
endmodule